`ifndef AXIS_TYPE_TEST_SVH
`define AXIS_TYPE_TEST_SVH

parameter DEST_WIDTH = 8;
parameter USER_WIDTH = 4;
parameter ID_WIDTH   = 4;

`include "axis_type.svh"

`endif
