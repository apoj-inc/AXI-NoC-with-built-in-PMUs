`define TEST

`include "axi_type_test.svh"
`include "axis_type_test.svh"
